library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity moving_average_tb is
end moving_average_tb;

architecture arch_moving_average_tb of moving_average_tb is
	
component moving_average is
generic (
  data_bits                     : integer := 8;
  group_length              : integer := 2 );
port (  i_clk                      : in  std_logic;
  -- input
  i_data                     : in  std_logic_vector(data_bits-1 downto 0);
  -- output
  --output the sum of group value
  o_data                     : out std_logic_vector(data_bits+group_length downto 0);
  oldest_data		     : out std_logic_vector(data_bits-1 downto 0));

end component moving_average;	
	

constant data_bits: integer := 8;
constant group_length: integer :=2;
signal  i_clk_tb:  std_logic:='0';
signal  i_data_tb: std_logic_vector(data_bits-1 downto 0):=(others=>'0');
signal  o_data_tb: std_logic_vector(data_bits+group_length downto 0):=(others=>'0');
signal  oldest_data_tb: std_logic_vector(data_bits-1 downto 0):=(others=>'0');
signal runsim : boolean := true;


begin
moving_average_component:

	component moving_average

	port map(
			i_clk =>i_clk_tb,
			i_data=>i_data_tb,
			o_data=>o_data_tb,
			oldest_data=>oldest_data_tb
);

    process
    begin
        if runsim then
            i_clk_tb <= '1';
            wait for 5 ns;
            i_clk_tb <= '0';
            wait for 5 ns;
        else
            wait;
        end if;
    end process;


test_process: process is
begin

wait for 13 ns;
i_data_tb <=x"01";
wait for 10 ns;
i_data_tb <=x"02";
wait for 10 ns;
i_data_tb <=x"03";
wait for 10 ns;
i_data_tb <=x"04";
wait for 10 ns;
i_data_tb <=x"05";
wait for 10 ns;
i_data_tb <=x"06";
wait for 10 ns;
i_data_tb <=x"07";
wait for 10 ns;
i_data_tb <=x"08";
wait for 10 ns;
i_data_tb <=x"09";
wait for 10 ns;
i_data_tb <=x"0A";

end process test_process;
end  arch_moving_average_tb;








